bind zad1 zad1_checker c0(.clk(clk), 
						  .rst(rst), 
						  .a(a), 
						  .b(b),  
						  .c(c), 
						  .d(d),  
						  .e(e), 
						  .f(f),  
						  .h(h), 
						  .g(g), 
						  .o1(o1), 
						  .o2(o2));
